// Copyright (C) 2018  Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License 
// Subscription Agreement, the Intel Quartus Prime License Agreement,
// the Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is for
// the sole purpose of programming logic devices manufactured by
// Intel and sold by Intel or its authorized distributors.  Please
// refer to the applicable agreement for further details.

// *****************************************************************************
// This file contains a Verilog test bench template that is freely editable to  
// suit user's needs .Comments are provided in each section to help the user    
// fill out necessary details.                                                  
// *****************************************************************************
// Generated on "10/05/2022 20:19:24"
                                                                                
// Verilog Test Bench template for design : phase_ramp_gen
// 
// Simulation tool : ModelSim-Altera (Verilog)
// 

`timescale 1 ns/ 100 ps
module phase_ramp_gen_tb();
// constants                                           
// general purpose registers
reg eachvec;
// test vector input registers
reg i_clk;
reg [31:0] i_fb_on;
reg [3:0] i_gain_sel;
reg [31:0] i_mod;
reg i_rst_n;
reg [31:0] i_step;
reg i_trig;
// wires                                               
wire o_change;
wire [31:0]  o_gain_sel2;
wire [31:0]  o_ladderWave;
wire [31:0]  o_phaseRamp;
wire [3:0]  o_shift_idx;
wire [1:0]  o_status;
wire [31:0]  o_step_init;

// assign statements (if any)                          
phase_ramp_gen i1 (
// port map - connection between master ports and signals/registers   
	.i_clk(i_clk),
	.i_fb_on(i_fb_on),
	.i_gain_sel(i_gain_sel),
	.i_mod(i_mod),
	.i_rst_n(i_rst_n),
	.i_step(i_step),
	.i_trig(i_trig),
	.o_change(o_change),
	.o_gain_sel2(o_gain_sel2),
	.o_ladderWave(o_ladderWave),
	.o_phaseRamp(o_phaseRamp),
	.o_shift_idx(o_shift_idx),
	.o_status(o_status),
	.o_step_init(o_step_init)
);
initial                                                
begin                                                  
// code that executes only once                        
// insert code here --> begin                          
                                                       
// --> end                                             
$display("Running testbench");                       
end                                                    
always                                                 
// optional sensitivity list                           
// @(event1 or event2 or .... eventn)                  
begin                                                  
// code executes for every event on sensitivity list   
// insert code here --> begin                          
                                                       
@eachvec;                                              
// --> end                                             
end                                                    
endmodule

