// CPU.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module CPU (
		input  wire        clk_clk,                  //      clk.clk
		output wire        dac_rst_export,           //  dac_rst.export
		output wire        epcs_dclk,                //     epcs.dclk
		output wire        epcs_sce,                 //         .sce
		output wire        epcs_sdo,                 //         .sdo
		input  wire        epcs_data0,               //         .data0
		input  wire        reset_reset_n,            //    reset.reset_n
		output wire [11:0] sdram_addr,               //    sdram.addr
		output wire [1:0]  sdram_ba,                 //         .ba
		output wire        sdram_cas_n,              //         .cas_n
		output wire        sdram_cke,                //         .cke
		output wire        sdram_cs_n,               //         .cs_n
		inout  wire [15:0] sdram_dq,                 //         .dq
		output wire [1:0]  sdram_dqm,                //         .dqm
		output wire        sdram_ras_n,              //         .ras_n
		output wire        sdram_we_n,               //         .we_n
		input  wire        spi_adc_MISO,             //  spi_adc.MISO
		output wire        spi_adc_MOSI,             //         .MOSI
		output wire        spi_adc_SCLK,             //         .SCLK
		output wire        spi_adc_SS_n,             //         .SS_n
		input  wire        spi_dac_MISO,             //  spi_dac.MISO
		output wire        spi_dac_MOSI,             //         .MOSI
		output wire        spi_dac_SCLK,             //         .SCLK
		output wire        spi_dac_SS_n,             //         .SS_n
		input  wire        sync_in_export,           //  sync_in.export
		input  wire        uart_rxd,                 //     uart.rxd
		output wire        uart_txd,                 //         .txd
		input  wire        uart_dbg_rxd,             // uart_dbg.rxd
		output wire        uart_dbg_txd,             //         .txd
		input  wire [31:0] varset_1_i_var0,          // varset_1.i_var0
		input  wire [31:0] varset_1_i_var1,          //         .i_var1
		input  wire [31:0] varset_1_i_var2,          //         .i_var2
		input  wire [31:0] varset_1_i_var3,          //         .i_var3
		input  wire [31:0] varset_1_i_var4,          //         .i_var4
		input  wire [31:0] varset_1_i_var5,          //         .i_var5
		input  wire [31:0] varset_1_i_var6,          //         .i_var6
		input  wire [31:0] varset_1_i_var7,          //         .i_var7
		input  wire [31:0] varset_1_i_var8,          //         .i_var8
		input  wire [31:0] varset_1_i_var9,          //         .i_var9
		input  wire [31:0] varset_1_i_var10,         //         .i_var10
		input  wire [31:0] varset_1_i_var11,         //         .i_var11
		input  wire [31:0] varset_1_i_var12,         //         .i_var12
		input  wire [31:0] varset_1_i_var13,         //         .i_var13
		input  wire [31:0] varset_1_i_var14,         //         .i_var14
		input  wire [31:0] varset_1_i_var15,         //         .i_var15
		input  wire [31:0] varset_1_i_var16,         //         .i_var16
		input  wire [31:0] varset_1_i_var17,         //         .i_var17
		input  wire [31:0] varset_1_i_var18,         //         .i_var18
		input  wire [31:0] varset_1_i_var19,         //         .i_var19
		input  wire [31:0] varset_1_i_var20,         //         .i_var20
		input  wire [31:0] varset_1_i_var21,         //         .i_var21
		input  wire [31:0] varset_1_i_var22,         //         .i_var22
		input  wire [31:0] varset_1_i_var23,         //         .i_var23
		input  wire [31:0] varset_1_i_var24,         //         .i_var24
		input  wire [31:0] varset_1_i_var25,         //         .i_var25
		input  wire [31:0] varset_1_i_var26,         //         .i_var26
		input  wire [31:0] varset_1_i_var27,         //         .i_var27
		input  wire [31:0] varset_1_i_var28,         //         .i_var28
		input  wire [31:0] varset_1_i_var29,         //         .i_var29
		input  wire [31:0] varset_1_i_var30,         //         .i_var30
		input  wire [31:0] varset_1_i_var31,         //         .i_var31
		input  wire [31:0] varset_1_i_var32,         //         .i_var32
		input  wire [31:0] varset_1_i_var33,         //         .i_var33
		input  wire [31:0] varset_1_i_var34,         //         .i_var34
		input  wire [31:0] varset_1_i_var35,         //         .i_var35
		input  wire [31:0] varset_1_i_var36,         //         .i_var36
		input  wire [31:0] varset_1_i_var37,         //         .i_var37
		input  wire [31:0] varset_1_i_var38,         //         .i_var38
		input  wire [31:0] varset_1_i_var39,         //         .i_var39
		input  wire [31:0] varset_1_i_var40,         //         .i_var40
		input  wire [31:0] varset_1_i_var41,         //         .i_var41
		input  wire [31:0] varset_1_i_var42,         //         .i_var42
		input  wire [31:0] varset_1_i_var43,         //         .i_var43
		input  wire [31:0] varset_1_i_var44,         //         .i_var44
		input  wire [31:0] varset_1_i_var45,         //         .i_var45
		input  wire [31:0] varset_1_i_var46,         //         .i_var46
		input  wire [31:0] varset_1_i_var47,         //         .i_var47
		input  wire [31:0] varset_1_i_var48,         //         .i_var48
		input  wire [31:0] varset_1_i_var49,         //         .i_var49
		input  wire [31:0] varset_1_i_var50,         //         .i_var50
		input  wire [31:0] varset_1_i_var51,         //         .i_var51
		input  wire [31:0] varset_1_i_var52,         //         .i_var52
		input  wire [31:0] varset_1_i_var53,         //         .i_var53
		input  wire [31:0] varset_1_i_var54,         //         .i_var54
		input  wire [31:0] varset_1_i_var55,         //         .i_var55
		input  wire [31:0] varset_1_i_var56,         //         .i_var56
		input  wire [31:0] varset_1_i_var57,         //         .i_var57
		input  wire [31:0] varset_1_i_var58,         //         .i_var58
		input  wire [31:0] varset_1_i_var59,         //         .i_var59
		output wire [31:0] varset_1_o_reg0,          //         .o_reg0
		output wire [31:0] varset_1_o_reg1,          //         .o_reg1
		output wire [31:0] varset_1_o_reg2,          //         .o_reg2
		output wire [31:0] varset_1_o_reg3,          //         .o_reg3
		output wire [31:0] varset_1_o_reg4,          //         .o_reg4
		output wire [31:0] varset_1_o_reg5,          //         .o_reg5
		output wire [31:0] varset_1_o_reg6,          //         .o_reg6
		output wire [31:0] varset_1_o_reg7,          //         .o_reg7
		output wire [31:0] varset_1_o_reg8,          //         .o_reg8
		output wire [31:0] varset_1_o_reg9,          //         .o_reg9
		output wire [31:0] varset_1_o_reg10,         //         .o_reg10
		output wire [31:0] varset_1_o_reg11,         //         .o_reg11
		output wire [31:0] varset_1_o_reg12,         //         .o_reg12
		output wire [31:0] varset_1_o_reg13,         //         .o_reg13
		output wire [31:0] varset_1_o_reg14,         //         .o_reg14
		output wire [31:0] varset_1_o_reg15,         //         .o_reg15
		output wire [31:0] varset_1_o_reg16,         //         .o_reg16
		output wire [31:0] varset_1_o_reg17,         //         .o_reg17
		output wire [31:0] varset_1_o_reg18,         //         .o_reg18
		output wire [31:0] varset_1_o_reg19,         //         .o_reg19
		output wire [31:0] varset_1_o_reg20,         //         .o_reg20
		output wire [31:0] varset_1_o_reg21,         //         .o_reg21
		output wire [31:0] varset_1_o_reg22,         //         .o_reg22
		output wire [31:0] varset_1_o_reg23,         //         .o_reg23
		output wire [31:0] varset_1_o_reg24,         //         .o_reg24
		output wire [31:0] varset_1_o_reg25,         //         .o_reg25
		output wire [31:0] varset_1_o_reg26,         //         .o_reg26
		output wire [31:0] varset_1_o_reg27,         //         .o_reg27
		output wire [31:0] varset_1_o_reg28,         //         .o_reg28
		output wire [31:0] varset_1_o_reg29,         //         .o_reg29
		output wire [31:0] varset_1_o_reg30,         //         .o_reg30
		output wire [31:0] varset_1_o_reg31,         //         .o_reg31
		output wire [31:0] varset_1_o_reg32,         //         .o_reg32
		output wire [31:0] varset_1_o_reg33,         //         .o_reg33
		output wire [31:0] varset_1_o_reg34,         //         .o_reg34
		output wire [31:0] varset_1_o_reg35,         //         .o_reg35
		output wire [31:0] varset_1_o_reg36,         //         .o_reg36
		output wire [31:0] varset_1_o_reg37,         //         .o_reg37
		output wire [31:0] varset_1_o_reg38,         //         .o_reg38
		output wire [31:0] varset_1_o_reg39,         //         .o_reg39
		output wire [31:0] varset_1_o_reg40,         //         .o_reg40
		output wire [31:0] varset_1_o_reg41,         //         .o_reg41
		output wire [31:0] varset_1_o_reg42,         //         .o_reg42
		output wire [31:0] varset_1_o_reg43,         //         .o_reg43
		output wire [31:0] varset_1_o_reg44,         //         .o_reg44
		output wire [31:0] varset_1_o_reg45,         //         .o_reg45
		output wire [31:0] varset_1_o_reg46,         //         .o_reg46
		output wire [31:0] varset_1_o_reg47,         //         .o_reg47
		output wire [31:0] varset_1_o_reg48,         //         .o_reg48
		output wire [31:0] varset_1_o_reg49,         //         .o_reg49
		output wire [31:0] varset_1_o_reg50,         //         .o_reg50
		output wire [31:0] varset_1_o_reg51,         //         .o_reg51
		output wire [31:0] varset_1_o_reg52,         //         .o_reg52
		output wire [31:0] varset_1_o_reg53,         //         .o_reg53
		output wire [31:0] varset_1_o_reg54,         //         .o_reg54
		output wire [31:0] varset_1_o_reg55,         //         .o_reg55
		output wire [31:0] varset_1_o_reg56,         //         .o_reg56
		output wire [31:0] varset_1_o_reg57,         //         .o_reg57
		output wire [31:0] varset_1_o_reg58,         //         .o_reg58
		output wire [31:0] varset_1_o_reg59,         //         .o_reg59
		output wire        varset_1_o_latch_trigger  //         .o_latch_trigger
	);

	wire  [31:0] nios2_data_master_readdata;                                // mm_interconnect_0:nios2_data_master_readdata -> nios2:d_readdata
	wire         nios2_data_master_waitrequest;                             // mm_interconnect_0:nios2_data_master_waitrequest -> nios2:d_waitrequest
	wire         nios2_data_master_debugaccess;                             // nios2:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_data_master_debugaccess
	wire  [25:0] nios2_data_master_address;                                 // nios2:d_address -> mm_interconnect_0:nios2_data_master_address
	wire   [3:0] nios2_data_master_byteenable;                              // nios2:d_byteenable -> mm_interconnect_0:nios2_data_master_byteenable
	wire         nios2_data_master_read;                                    // nios2:d_read -> mm_interconnect_0:nios2_data_master_read
	wire         nios2_data_master_write;                                   // nios2:d_write -> mm_interconnect_0:nios2_data_master_write
	wire  [31:0] nios2_data_master_writedata;                               // nios2:d_writedata -> mm_interconnect_0:nios2_data_master_writedata
	wire  [31:0] nios2_instruction_master_readdata;                         // mm_interconnect_0:nios2_instruction_master_readdata -> nios2:i_readdata
	wire         nios2_instruction_master_waitrequest;                      // mm_interconnect_0:nios2_instruction_master_waitrequest -> nios2:i_waitrequest
	wire  [25:0] nios2_instruction_master_address;                          // nios2:i_address -> mm_interconnect_0:nios2_instruction_master_address
	wire         nios2_instruction_master_read;                             // nios2:i_read -> mm_interconnect_0:nios2_instruction_master_read
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;    // jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest; // jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire         mm_interconnect_0_varset_1_avalon_slave_chipselect;        // mm_interconnect_0:VarSet_1_avalon_slave_chipselect -> VarSet_1:chipselect
	wire  [31:0] mm_interconnect_0_varset_1_avalon_slave_readdata;          // VarSet_1:readdata -> mm_interconnect_0:VarSet_1_avalon_slave_readdata
	wire   [6:0] mm_interconnect_0_varset_1_avalon_slave_address;           // mm_interconnect_0:VarSet_1_avalon_slave_address -> VarSet_1:address
	wire         mm_interconnect_0_varset_1_avalon_slave_write;             // mm_interconnect_0:VarSet_1_avalon_slave_write -> VarSet_1:write_n
	wire  [31:0] mm_interconnect_0_varset_1_avalon_slave_writedata;         // mm_interconnect_0:VarSet_1_avalon_slave_writedata -> VarSet_1:writedata
	wire  [31:0] mm_interconnect_0_sysid_control_slave_readdata;            // sysid:readdata -> mm_interconnect_0:sysid_control_slave_readdata
	wire   [0:0] mm_interconnect_0_sysid_control_slave_address;             // mm_interconnect_0:sysid_control_slave_address -> sysid:address
	wire  [31:0] mm_interconnect_0_nios2_debug_mem_slave_readdata;          // nios2:debug_mem_slave_readdata -> mm_interconnect_0:nios2_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios2_debug_mem_slave_waitrequest;       // nios2:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios2_debug_mem_slave_debugaccess;       // mm_interconnect_0:nios2_debug_mem_slave_debugaccess -> nios2:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_debug_mem_slave_address;           // mm_interconnect_0:nios2_debug_mem_slave_address -> nios2:debug_mem_slave_address
	wire         mm_interconnect_0_nios2_debug_mem_slave_read;              // mm_interconnect_0:nios2_debug_mem_slave_read -> nios2:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios2_debug_mem_slave_byteenable;        // mm_interconnect_0:nios2_debug_mem_slave_byteenable -> nios2:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios2_debug_mem_slave_write;             // mm_interconnect_0:nios2_debug_mem_slave_write -> nios2:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios2_debug_mem_slave_writedata;         // mm_interconnect_0:nios2_debug_mem_slave_writedata -> nios2:debug_mem_slave_writedata
	wire         mm_interconnect_0_epcs_epcs_control_port_chipselect;       // mm_interconnect_0:epcs_epcs_control_port_chipselect -> epcs:chipselect
	wire  [31:0] mm_interconnect_0_epcs_epcs_control_port_readdata;         // epcs:readdata -> mm_interconnect_0:epcs_epcs_control_port_readdata
	wire   [8:0] mm_interconnect_0_epcs_epcs_control_port_address;          // mm_interconnect_0:epcs_epcs_control_port_address -> epcs:address
	wire         mm_interconnect_0_epcs_epcs_control_port_read;             // mm_interconnect_0:epcs_epcs_control_port_read -> epcs:read_n
	wire         mm_interconnect_0_epcs_epcs_control_port_write;            // mm_interconnect_0:epcs_epcs_control_port_write -> epcs:write_n
	wire  [31:0] mm_interconnect_0_epcs_epcs_control_port_writedata;        // mm_interconnect_0:epcs_epcs_control_port_writedata -> epcs:writedata
	wire         mm_interconnect_0_sdram_s1_chipselect;                     // mm_interconnect_0:sdram_s1_chipselect -> sdram:az_cs
	wire  [15:0] mm_interconnect_0_sdram_s1_readdata;                       // sdram:za_data -> mm_interconnect_0:sdram_s1_readdata
	wire         mm_interconnect_0_sdram_s1_waitrequest;                    // sdram:za_waitrequest -> mm_interconnect_0:sdram_s1_waitrequest
	wire  [22:0] mm_interconnect_0_sdram_s1_address;                        // mm_interconnect_0:sdram_s1_address -> sdram:az_addr
	wire         mm_interconnect_0_sdram_s1_read;                           // mm_interconnect_0:sdram_s1_read -> sdram:az_rd_n
	wire   [1:0] mm_interconnect_0_sdram_s1_byteenable;                     // mm_interconnect_0:sdram_s1_byteenable -> sdram:az_be_n
	wire         mm_interconnect_0_sdram_s1_readdatavalid;                  // sdram:za_valid -> mm_interconnect_0:sdram_s1_readdatavalid
	wire         mm_interconnect_0_sdram_s1_write;                          // mm_interconnect_0:sdram_s1_write -> sdram:az_wr_n
	wire  [15:0] mm_interconnect_0_sdram_s1_writedata;                      // mm_interconnect_0:sdram_s1_writedata -> sdram:az_data
	wire         mm_interconnect_0_sync_in_s1_chipselect;                   // mm_interconnect_0:sync_in_s1_chipselect -> sync_in:chipselect
	wire  [31:0] mm_interconnect_0_sync_in_s1_readdata;                     // sync_in:readdata -> mm_interconnect_0:sync_in_s1_readdata
	wire   [1:0] mm_interconnect_0_sync_in_s1_address;                      // mm_interconnect_0:sync_in_s1_address -> sync_in:address
	wire         mm_interconnect_0_sync_in_s1_write;                        // mm_interconnect_0:sync_in_s1_write -> sync_in:write_n
	wire  [31:0] mm_interconnect_0_sync_in_s1_writedata;                    // mm_interconnect_0:sync_in_s1_writedata -> sync_in:writedata
	wire         mm_interconnect_0_uart_s1_chipselect;                      // mm_interconnect_0:uart_s1_chipselect -> uart:chipselect
	wire  [15:0] mm_interconnect_0_uart_s1_readdata;                        // uart:readdata -> mm_interconnect_0:uart_s1_readdata
	wire   [2:0] mm_interconnect_0_uart_s1_address;                         // mm_interconnect_0:uart_s1_address -> uart:address
	wire         mm_interconnect_0_uart_s1_read;                            // mm_interconnect_0:uart_s1_read -> uart:read_n
	wire         mm_interconnect_0_uart_s1_begintransfer;                   // mm_interconnect_0:uart_s1_begintransfer -> uart:begintransfer
	wire         mm_interconnect_0_uart_s1_write;                           // mm_interconnect_0:uart_s1_write -> uart:write_n
	wire  [15:0] mm_interconnect_0_uart_s1_writedata;                       // mm_interconnect_0:uart_s1_writedata -> uart:writedata
	wire         mm_interconnect_0_uart_dbg_s1_chipselect;                  // mm_interconnect_0:uart_dbg_s1_chipselect -> uart_dbg:chipselect
	wire  [15:0] mm_interconnect_0_uart_dbg_s1_readdata;                    // uart_dbg:readdata -> mm_interconnect_0:uart_dbg_s1_readdata
	wire   [2:0] mm_interconnect_0_uart_dbg_s1_address;                     // mm_interconnect_0:uart_dbg_s1_address -> uart_dbg:address
	wire         mm_interconnect_0_uart_dbg_s1_read;                        // mm_interconnect_0:uart_dbg_s1_read -> uart_dbg:read_n
	wire         mm_interconnect_0_uart_dbg_s1_begintransfer;               // mm_interconnect_0:uart_dbg_s1_begintransfer -> uart_dbg:begintransfer
	wire         mm_interconnect_0_uart_dbg_s1_write;                       // mm_interconnect_0:uart_dbg_s1_write -> uart_dbg:write_n
	wire  [15:0] mm_interconnect_0_uart_dbg_s1_writedata;                   // mm_interconnect_0:uart_dbg_s1_writedata -> uart_dbg:writedata
	wire         mm_interconnect_0_dac_rst_s1_chipselect;                   // mm_interconnect_0:DAC_RST_s1_chipselect -> DAC_RST:chipselect
	wire  [31:0] mm_interconnect_0_dac_rst_s1_readdata;                     // DAC_RST:readdata -> mm_interconnect_0:DAC_RST_s1_readdata
	wire   [1:0] mm_interconnect_0_dac_rst_s1_address;                      // mm_interconnect_0:DAC_RST_s1_address -> DAC_RST:address
	wire         mm_interconnect_0_dac_rst_s1_write;                        // mm_interconnect_0:DAC_RST_s1_write -> DAC_RST:write_n
	wire  [31:0] mm_interconnect_0_dac_rst_s1_writedata;                    // mm_interconnect_0:DAC_RST_s1_writedata -> DAC_RST:writedata
	wire         mm_interconnect_0_spi_adc_spi_control_port_chipselect;     // mm_interconnect_0:spi_ADC_spi_control_port_chipselect -> spi_ADC:spi_select
	wire  [15:0] mm_interconnect_0_spi_adc_spi_control_port_readdata;       // spi_ADC:data_to_cpu -> mm_interconnect_0:spi_ADC_spi_control_port_readdata
	wire   [2:0] mm_interconnect_0_spi_adc_spi_control_port_address;        // mm_interconnect_0:spi_ADC_spi_control_port_address -> spi_ADC:mem_addr
	wire         mm_interconnect_0_spi_adc_spi_control_port_read;           // mm_interconnect_0:spi_ADC_spi_control_port_read -> spi_ADC:read_n
	wire         mm_interconnect_0_spi_adc_spi_control_port_write;          // mm_interconnect_0:spi_ADC_spi_control_port_write -> spi_ADC:write_n
	wire  [15:0] mm_interconnect_0_spi_adc_spi_control_port_writedata;      // mm_interconnect_0:spi_ADC_spi_control_port_writedata -> spi_ADC:data_from_cpu
	wire         mm_interconnect_0_spi_dac_spi_control_port_chipselect;     // mm_interconnect_0:spi_DAC_spi_control_port_chipselect -> spi_DAC:spi_select
	wire  [15:0] mm_interconnect_0_spi_dac_spi_control_port_readdata;       // spi_DAC:data_to_cpu -> mm_interconnect_0:spi_DAC_spi_control_port_readdata
	wire   [2:0] mm_interconnect_0_spi_dac_spi_control_port_address;        // mm_interconnect_0:spi_DAC_spi_control_port_address -> spi_DAC:mem_addr
	wire         mm_interconnect_0_spi_dac_spi_control_port_read;           // mm_interconnect_0:spi_DAC_spi_control_port_read -> spi_DAC:read_n
	wire         mm_interconnect_0_spi_dac_spi_control_port_write;          // mm_interconnect_0:spi_DAC_spi_control_port_write -> spi_DAC:write_n
	wire  [15:0] mm_interconnect_0_spi_dac_spi_control_port_writedata;      // mm_interconnect_0:spi_DAC_spi_control_port_writedata -> spi_DAC:data_from_cpu
	wire         irq_mapper_receiver0_irq;                                  // jtag_uart:av_irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                  // spi_ADC:irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                  // epcs:irq -> irq_mapper:receiver2_irq
	wire         irq_mapper_receiver3_irq;                                  // sync_in:irq -> irq_mapper:receiver3_irq
	wire         irq_mapper_receiver4_irq;                                  // uart:irq -> irq_mapper:receiver4_irq
	wire         irq_mapper_receiver5_irq;                                  // uart_dbg:irq -> irq_mapper:receiver5_irq
	wire         irq_mapper_receiver6_irq;                                  // spi_DAC:irq -> irq_mapper:receiver6_irq
	wire  [31:0] nios2_irq_irq;                                             // irq_mapper:sender_irq -> nios2:irq
	wire         rst_controller_reset_out_reset;                            // rst_controller:reset_out -> [DAC_RST:reset_n, VarSet_1:rst_n, epcs:reset_n, mm_interconnect_0:VarSet_1_reset_n_reset_bridge_in_reset_reset, rst_translator:in_reset, sdram:reset_n, spi_ADC:reset_n, spi_DAC:reset_n, sync_in:reset_n, sysid:reset_n, uart:reset_n, uart_dbg:reset_n]
	wire         rst_controller_reset_out_reset_req;                        // rst_controller:reset_req -> [epcs:reset_req, rst_translator:reset_req_in]
	wire         nios2_debug_reset_request_reset;                           // nios2:debug_reset_request -> rst_controller:reset_in1
	wire         rst_controller_001_reset_out_reset;                        // rst_controller_001:reset_out -> [irq_mapper:reset, jtag_uart:rst_n, mm_interconnect_0:nios2_reset_reset_bridge_in_reset_reset, nios2:reset_n, rst_translator_001:in_reset]
	wire         rst_controller_001_reset_out_reset_req;                    // rst_controller_001:reset_req -> [nios2:reset_req, rst_translator_001:reset_req_in]

	CPU_DAC_RST dac_rst (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_dac_rst_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_dac_rst_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_dac_rst_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_dac_rst_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_dac_rst_s1_readdata),   //                    .readdata
		.out_port   (dac_rst_export)                           // external_connection.export
	);

	GyroVarSet_60 varset_1 (
		.clk             (clk_clk),                                            //        clock.clk
		.rst_n           (~rst_controller_reset_out_reset),                    //      reset_n.reset_n
		.address         (mm_interconnect_0_varset_1_avalon_slave_address),    // avalon_slave.address
		.chipselect      (mm_interconnect_0_varset_1_avalon_slave_chipselect), //             .chipselect
		.write_n         (~mm_interconnect_0_varset_1_avalon_slave_write),     //             .write_n
		.writedata       (mm_interconnect_0_varset_1_avalon_slave_writedata),  //             .writedata
		.readdata        (mm_interconnect_0_varset_1_avalon_slave_readdata),   //             .readdata
		.i_var0          (varset_1_i_var0),                                    //      conduit.i_var0
		.i_var1          (varset_1_i_var1),                                    //             .i_var1
		.i_var2          (varset_1_i_var2),                                    //             .i_var2
		.i_var3          (varset_1_i_var3),                                    //             .i_var3
		.i_var4          (varset_1_i_var4),                                    //             .i_var4
		.i_var5          (varset_1_i_var5),                                    //             .i_var5
		.i_var6          (varset_1_i_var6),                                    //             .i_var6
		.i_var7          (varset_1_i_var7),                                    //             .i_var7
		.i_var8          (varset_1_i_var8),                                    //             .i_var8
		.i_var9          (varset_1_i_var9),                                    //             .i_var9
		.i_var10         (varset_1_i_var10),                                   //             .i_var10
		.i_var11         (varset_1_i_var11),                                   //             .i_var11
		.i_var12         (varset_1_i_var12),                                   //             .i_var12
		.i_var13         (varset_1_i_var13),                                   //             .i_var13
		.i_var14         (varset_1_i_var14),                                   //             .i_var14
		.i_var15         (varset_1_i_var15),                                   //             .i_var15
		.i_var16         (varset_1_i_var16),                                   //             .i_var16
		.i_var17         (varset_1_i_var17),                                   //             .i_var17
		.i_var18         (varset_1_i_var18),                                   //             .i_var18
		.i_var19         (varset_1_i_var19),                                   //             .i_var19
		.i_var20         (varset_1_i_var20),                                   //             .i_var20
		.i_var21         (varset_1_i_var21),                                   //             .i_var21
		.i_var22         (varset_1_i_var22),                                   //             .i_var22
		.i_var23         (varset_1_i_var23),                                   //             .i_var23
		.i_var24         (varset_1_i_var24),                                   //             .i_var24
		.i_var25         (varset_1_i_var25),                                   //             .i_var25
		.i_var26         (varset_1_i_var26),                                   //             .i_var26
		.i_var27         (varset_1_i_var27),                                   //             .i_var27
		.i_var28         (varset_1_i_var28),                                   //             .i_var28
		.i_var29         (varset_1_i_var29),                                   //             .i_var29
		.i_var30         (varset_1_i_var30),                                   //             .i_var30
		.i_var31         (varset_1_i_var31),                                   //             .i_var31
		.i_var32         (varset_1_i_var32),                                   //             .i_var32
		.i_var33         (varset_1_i_var33),                                   //             .i_var33
		.i_var34         (varset_1_i_var34),                                   //             .i_var34
		.i_var35         (varset_1_i_var35),                                   //             .i_var35
		.i_var36         (varset_1_i_var36),                                   //             .i_var36
		.i_var37         (varset_1_i_var37),                                   //             .i_var37
		.i_var38         (varset_1_i_var38),                                   //             .i_var38
		.i_var39         (varset_1_i_var39),                                   //             .i_var39
		.i_var40         (varset_1_i_var40),                                   //             .i_var40
		.i_var41         (varset_1_i_var41),                                   //             .i_var41
		.i_var42         (varset_1_i_var42),                                   //             .i_var42
		.i_var43         (varset_1_i_var43),                                   //             .i_var43
		.i_var44         (varset_1_i_var44),                                   //             .i_var44
		.i_var45         (varset_1_i_var45),                                   //             .i_var45
		.i_var46         (varset_1_i_var46),                                   //             .i_var46
		.i_var47         (varset_1_i_var47),                                   //             .i_var47
		.i_var48         (varset_1_i_var48),                                   //             .i_var48
		.i_var49         (varset_1_i_var49),                                   //             .i_var49
		.i_var50         (varset_1_i_var50),                                   //             .i_var50
		.i_var51         (varset_1_i_var51),                                   //             .i_var51
		.i_var52         (varset_1_i_var52),                                   //             .i_var52
		.i_var53         (varset_1_i_var53),                                   //             .i_var53
		.i_var54         (varset_1_i_var54),                                   //             .i_var54
		.i_var55         (varset_1_i_var55),                                   //             .i_var55
		.i_var56         (varset_1_i_var56),                                   //             .i_var56
		.i_var57         (varset_1_i_var57),                                   //             .i_var57
		.i_var58         (varset_1_i_var58),                                   //             .i_var58
		.i_var59         (varset_1_i_var59),                                   //             .i_var59
		.o_reg0          (varset_1_o_reg0),                                    //             .o_reg0
		.o_reg1          (varset_1_o_reg1),                                    //             .o_reg1
		.o_reg2          (varset_1_o_reg2),                                    //             .o_reg2
		.o_reg3          (varset_1_o_reg3),                                    //             .o_reg3
		.o_reg4          (varset_1_o_reg4),                                    //             .o_reg4
		.o_reg5          (varset_1_o_reg5),                                    //             .o_reg5
		.o_reg6          (varset_1_o_reg6),                                    //             .o_reg6
		.o_reg7          (varset_1_o_reg7),                                    //             .o_reg7
		.o_reg8          (varset_1_o_reg8),                                    //             .o_reg8
		.o_reg9          (varset_1_o_reg9),                                    //             .o_reg9
		.o_reg10         (varset_1_o_reg10),                                   //             .o_reg10
		.o_reg11         (varset_1_o_reg11),                                   //             .o_reg11
		.o_reg12         (varset_1_o_reg12),                                   //             .o_reg12
		.o_reg13         (varset_1_o_reg13),                                   //             .o_reg13
		.o_reg14         (varset_1_o_reg14),                                   //             .o_reg14
		.o_reg15         (varset_1_o_reg15),                                   //             .o_reg15
		.o_reg16         (varset_1_o_reg16),                                   //             .o_reg16
		.o_reg17         (varset_1_o_reg17),                                   //             .o_reg17
		.o_reg18         (varset_1_o_reg18),                                   //             .o_reg18
		.o_reg19         (varset_1_o_reg19),                                   //             .o_reg19
		.o_reg20         (varset_1_o_reg20),                                   //             .o_reg20
		.o_reg21         (varset_1_o_reg21),                                   //             .o_reg21
		.o_reg22         (varset_1_o_reg22),                                   //             .o_reg22
		.o_reg23         (varset_1_o_reg23),                                   //             .o_reg23
		.o_reg24         (varset_1_o_reg24),                                   //             .o_reg24
		.o_reg25         (varset_1_o_reg25),                                   //             .o_reg25
		.o_reg26         (varset_1_o_reg26),                                   //             .o_reg26
		.o_reg27         (varset_1_o_reg27),                                   //             .o_reg27
		.o_reg28         (varset_1_o_reg28),                                   //             .o_reg28
		.o_reg29         (varset_1_o_reg29),                                   //             .o_reg29
		.o_reg30         (varset_1_o_reg30),                                   //             .o_reg30
		.o_reg31         (varset_1_o_reg31),                                   //             .o_reg31
		.o_reg32         (varset_1_o_reg32),                                   //             .o_reg32
		.o_reg33         (varset_1_o_reg33),                                   //             .o_reg33
		.o_reg34         (varset_1_o_reg34),                                   //             .o_reg34
		.o_reg35         (varset_1_o_reg35),                                   //             .o_reg35
		.o_reg36         (varset_1_o_reg36),                                   //             .o_reg36
		.o_reg37         (varset_1_o_reg37),                                   //             .o_reg37
		.o_reg38         (varset_1_o_reg38),                                   //             .o_reg38
		.o_reg39         (varset_1_o_reg39),                                   //             .o_reg39
		.o_reg40         (varset_1_o_reg40),                                   //             .o_reg40
		.o_reg41         (varset_1_o_reg41),                                   //             .o_reg41
		.o_reg42         (varset_1_o_reg42),                                   //             .o_reg42
		.o_reg43         (varset_1_o_reg43),                                   //             .o_reg43
		.o_reg44         (varset_1_o_reg44),                                   //             .o_reg44
		.o_reg45         (varset_1_o_reg45),                                   //             .o_reg45
		.o_reg46         (varset_1_o_reg46),                                   //             .o_reg46
		.o_reg47         (varset_1_o_reg47),                                   //             .o_reg47
		.o_reg48         (varset_1_o_reg48),                                   //             .o_reg48
		.o_reg49         (varset_1_o_reg49),                                   //             .o_reg49
		.o_reg50         (varset_1_o_reg50),                                   //             .o_reg50
		.o_reg51         (varset_1_o_reg51),                                   //             .o_reg51
		.o_reg52         (varset_1_o_reg52),                                   //             .o_reg52
		.o_reg53         (varset_1_o_reg53),                                   //             .o_reg53
		.o_reg54         (varset_1_o_reg54),                                   //             .o_reg54
		.o_reg55         (varset_1_o_reg55),                                   //             .o_reg55
		.o_reg56         (varset_1_o_reg56),                                   //             .o_reg56
		.o_reg57         (varset_1_o_reg57),                                   //             .o_reg57
		.o_reg58         (varset_1_o_reg58),                                   //             .o_reg58
		.o_reg59         (varset_1_o_reg59),                                   //             .o_reg59
		.o_latch_trigger (varset_1_o_latch_trigger)                            //             .o_latch_trigger
	);

	CPU_epcs epcs (
		.clk        (clk_clk),                                             //               clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                     //             reset.reset_n
		.reset_req  (rst_controller_reset_out_reset_req),                  //                  .reset_req
		.address    (mm_interconnect_0_epcs_epcs_control_port_address),    // epcs_control_port.address
		.chipselect (mm_interconnect_0_epcs_epcs_control_port_chipselect), //                  .chipselect
		.read_n     (~mm_interconnect_0_epcs_epcs_control_port_read),      //                  .read_n
		.readdata   (mm_interconnect_0_epcs_epcs_control_port_readdata),   //                  .readdata
		.write_n    (~mm_interconnect_0_epcs_epcs_control_port_write),     //                  .write_n
		.writedata  (mm_interconnect_0_epcs_epcs_control_port_writedata),  //                  .writedata
		.irq        (irq_mapper_receiver2_irq),                            //               irq.irq
		.dclk       (epcs_dclk),                                           //          external.export
		.sce        (epcs_sce),                                            //                  .export
		.sdo        (epcs_sdo),                                            //                  .export
		.data0      (epcs_data0)                                           //                  .export
	);

	CPU_jtag_uart jtag_uart (
		.clk            (clk_clk),                                                   //               clk.clk
		.rst_n          (~rst_controller_001_reset_out_reset),                       //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                   //               irq.irq
	);

	CPU_nios2 nios2 (
		.clk                                 (clk_clk),                                             //                       clk.clk
		.reset_n                             (~rst_controller_001_reset_out_reset),                 //                     reset.reset_n
		.reset_req                           (rst_controller_001_reset_out_reset_req),              //                          .reset_req
		.d_address                           (nios2_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_data_master_read),                              //                          .read
		.d_readdata                          (nios2_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_data_master_write),                             //                          .write
		.d_writedata                         (nios2_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (nios2_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (nios2_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (nios2_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                     // custom_instruction_master.readra
	);

	CPU_sdram sdram (
		.clk            (clk_clk),                                  //   clk.clk
		.reset_n        (~rst_controller_reset_out_reset),          // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_addr),                               //  wire.export
		.zs_ba          (sdram_ba),                                 //      .export
		.zs_cas_n       (sdram_cas_n),                              //      .export
		.zs_cke         (sdram_cke),                                //      .export
		.zs_cs_n        (sdram_cs_n),                               //      .export
		.zs_dq          (sdram_dq),                                 //      .export
		.zs_dqm         (sdram_dqm),                                //      .export
		.zs_ras_n       (sdram_ras_n),                              //      .export
		.zs_we_n        (sdram_we_n)                                //      .export
	);

	CPU_spi_ADC spi_adc (
		.clk           (clk_clk),                                               //              clk.clk
		.reset_n       (~rst_controller_reset_out_reset),                       //            reset.reset_n
		.data_from_cpu (mm_interconnect_0_spi_adc_spi_control_port_writedata),  // spi_control_port.writedata
		.data_to_cpu   (mm_interconnect_0_spi_adc_spi_control_port_readdata),   //                 .readdata
		.mem_addr      (mm_interconnect_0_spi_adc_spi_control_port_address),    //                 .address
		.read_n        (~mm_interconnect_0_spi_adc_spi_control_port_read),      //                 .read_n
		.spi_select    (mm_interconnect_0_spi_adc_spi_control_port_chipselect), //                 .chipselect
		.write_n       (~mm_interconnect_0_spi_adc_spi_control_port_write),     //                 .write_n
		.irq           (irq_mapper_receiver1_irq),                              //              irq.irq
		.MISO          (spi_adc_MISO),                                          //         external.export
		.MOSI          (spi_adc_MOSI),                                          //                 .export
		.SCLK          (spi_adc_SCLK),                                          //                 .export
		.SS_n          (spi_adc_SS_n)                                           //                 .export
	);

	CPU_spi_ADC spi_dac (
		.clk           (clk_clk),                                               //              clk.clk
		.reset_n       (~rst_controller_reset_out_reset),                       //            reset.reset_n
		.data_from_cpu (mm_interconnect_0_spi_dac_spi_control_port_writedata),  // spi_control_port.writedata
		.data_to_cpu   (mm_interconnect_0_spi_dac_spi_control_port_readdata),   //                 .readdata
		.mem_addr      (mm_interconnect_0_spi_dac_spi_control_port_address),    //                 .address
		.read_n        (~mm_interconnect_0_spi_dac_spi_control_port_read),      //                 .read_n
		.spi_select    (mm_interconnect_0_spi_dac_spi_control_port_chipselect), //                 .chipselect
		.write_n       (~mm_interconnect_0_spi_dac_spi_control_port_write),     //                 .write_n
		.irq           (irq_mapper_receiver6_irq),                              //              irq.irq
		.MISO          (spi_dac_MISO),                                          //         external.export
		.MOSI          (spi_dac_MOSI),                                          //                 .export
		.SCLK          (spi_dac_SCLK),                                          //                 .export
		.SS_n          (spi_dac_SS_n)                                           //                 .export
	);

	CPU_sync_in sync_in (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_sync_in_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_sync_in_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_sync_in_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_sync_in_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_sync_in_s1_readdata),   //                    .readdata
		.in_port    (sync_in_export),                          // external_connection.export
		.irq        (irq_mapper_receiver3_irq)                 //                 irq.irq
	);

	CPU_sysid sysid (
		.clock    (clk_clk),                                        //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_control_slave_address)   //              .address
	);

	CPU_uart uart (
		.clk           (clk_clk),                                 //                 clk.clk
		.reset_n       (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address       (mm_interconnect_0_uart_s1_address),       //                  s1.address
		.begintransfer (mm_interconnect_0_uart_s1_begintransfer), //                    .begintransfer
		.chipselect    (mm_interconnect_0_uart_s1_chipselect),    //                    .chipselect
		.read_n        (~mm_interconnect_0_uart_s1_read),         //                    .read_n
		.write_n       (~mm_interconnect_0_uart_s1_write),        //                    .write_n
		.writedata     (mm_interconnect_0_uart_s1_writedata),     //                    .writedata
		.readdata      (mm_interconnect_0_uart_s1_readdata),      //                    .readdata
		.rxd           (uart_rxd),                                // external_connection.export
		.txd           (uart_txd),                                //                    .export
		.irq           (irq_mapper_receiver4_irq)                 //                 irq.irq
	);

	CPU_uart uart_dbg (
		.clk           (clk_clk),                                     //                 clk.clk
		.reset_n       (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address       (mm_interconnect_0_uart_dbg_s1_address),       //                  s1.address
		.begintransfer (mm_interconnect_0_uart_dbg_s1_begintransfer), //                    .begintransfer
		.chipselect    (mm_interconnect_0_uart_dbg_s1_chipselect),    //                    .chipselect
		.read_n        (~mm_interconnect_0_uart_dbg_s1_read),         //                    .read_n
		.write_n       (~mm_interconnect_0_uart_dbg_s1_write),        //                    .write_n
		.writedata     (mm_interconnect_0_uart_dbg_s1_writedata),     //                    .writedata
		.readdata      (mm_interconnect_0_uart_dbg_s1_readdata),      //                    .readdata
		.rxd           (uart_dbg_rxd),                                // external_connection.export
		.txd           (uart_dbg_txd),                                //                    .export
		.irq           (irq_mapper_receiver5_irq)                     //                 irq.irq
	);

	CPU_mm_interconnect_0 mm_interconnect_0 (
		.clk_CPU_clk_clk                              (clk_clk),                                                   //                            clk_CPU_clk.clk
		.nios2_reset_reset_bridge_in_reset_reset      (rst_controller_001_reset_out_reset),                        //      nios2_reset_reset_bridge_in_reset.reset
		.VarSet_1_reset_n_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                            // VarSet_1_reset_n_reset_bridge_in_reset.reset
		.nios2_data_master_address                    (nios2_data_master_address),                                 //                      nios2_data_master.address
		.nios2_data_master_waitrequest                (nios2_data_master_waitrequest),                             //                                       .waitrequest
		.nios2_data_master_byteenable                 (nios2_data_master_byteenable),                              //                                       .byteenable
		.nios2_data_master_read                       (nios2_data_master_read),                                    //                                       .read
		.nios2_data_master_readdata                   (nios2_data_master_readdata),                                //                                       .readdata
		.nios2_data_master_write                      (nios2_data_master_write),                                   //                                       .write
		.nios2_data_master_writedata                  (nios2_data_master_writedata),                               //                                       .writedata
		.nios2_data_master_debugaccess                (nios2_data_master_debugaccess),                             //                                       .debugaccess
		.nios2_instruction_master_address             (nios2_instruction_master_address),                          //               nios2_instruction_master.address
		.nios2_instruction_master_waitrequest         (nios2_instruction_master_waitrequest),                      //                                       .waitrequest
		.nios2_instruction_master_read                (nios2_instruction_master_read),                             //                                       .read
		.nios2_instruction_master_readdata            (nios2_instruction_master_readdata),                         //                                       .readdata
		.DAC_RST_s1_address                           (mm_interconnect_0_dac_rst_s1_address),                      //                             DAC_RST_s1.address
		.DAC_RST_s1_write                             (mm_interconnect_0_dac_rst_s1_write),                        //                                       .write
		.DAC_RST_s1_readdata                          (mm_interconnect_0_dac_rst_s1_readdata),                     //                                       .readdata
		.DAC_RST_s1_writedata                         (mm_interconnect_0_dac_rst_s1_writedata),                    //                                       .writedata
		.DAC_RST_s1_chipselect                        (mm_interconnect_0_dac_rst_s1_chipselect),                   //                                       .chipselect
		.epcs_epcs_control_port_address               (mm_interconnect_0_epcs_epcs_control_port_address),          //                 epcs_epcs_control_port.address
		.epcs_epcs_control_port_write                 (mm_interconnect_0_epcs_epcs_control_port_write),            //                                       .write
		.epcs_epcs_control_port_read                  (mm_interconnect_0_epcs_epcs_control_port_read),             //                                       .read
		.epcs_epcs_control_port_readdata              (mm_interconnect_0_epcs_epcs_control_port_readdata),         //                                       .readdata
		.epcs_epcs_control_port_writedata             (mm_interconnect_0_epcs_epcs_control_port_writedata),        //                                       .writedata
		.epcs_epcs_control_port_chipselect            (mm_interconnect_0_epcs_epcs_control_port_chipselect),       //                                       .chipselect
		.jtag_uart_avalon_jtag_slave_address          (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //            jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write            (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),       //                                       .write
		.jtag_uart_avalon_jtag_slave_read             (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),        //                                       .read
		.jtag_uart_avalon_jtag_slave_readdata         (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                                       .readdata
		.jtag_uart_avalon_jtag_slave_writedata        (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                                       .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest      (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                                       .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect       (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  //                                       .chipselect
		.nios2_debug_mem_slave_address                (mm_interconnect_0_nios2_debug_mem_slave_address),           //                  nios2_debug_mem_slave.address
		.nios2_debug_mem_slave_write                  (mm_interconnect_0_nios2_debug_mem_slave_write),             //                                       .write
		.nios2_debug_mem_slave_read                   (mm_interconnect_0_nios2_debug_mem_slave_read),              //                                       .read
		.nios2_debug_mem_slave_readdata               (mm_interconnect_0_nios2_debug_mem_slave_readdata),          //                                       .readdata
		.nios2_debug_mem_slave_writedata              (mm_interconnect_0_nios2_debug_mem_slave_writedata),         //                                       .writedata
		.nios2_debug_mem_slave_byteenable             (mm_interconnect_0_nios2_debug_mem_slave_byteenable),        //                                       .byteenable
		.nios2_debug_mem_slave_waitrequest            (mm_interconnect_0_nios2_debug_mem_slave_waitrequest),       //                                       .waitrequest
		.nios2_debug_mem_slave_debugaccess            (mm_interconnect_0_nios2_debug_mem_slave_debugaccess),       //                                       .debugaccess
		.sdram_s1_address                             (mm_interconnect_0_sdram_s1_address),                        //                               sdram_s1.address
		.sdram_s1_write                               (mm_interconnect_0_sdram_s1_write),                          //                                       .write
		.sdram_s1_read                                (mm_interconnect_0_sdram_s1_read),                           //                                       .read
		.sdram_s1_readdata                            (mm_interconnect_0_sdram_s1_readdata),                       //                                       .readdata
		.sdram_s1_writedata                           (mm_interconnect_0_sdram_s1_writedata),                      //                                       .writedata
		.sdram_s1_byteenable                          (mm_interconnect_0_sdram_s1_byteenable),                     //                                       .byteenable
		.sdram_s1_readdatavalid                       (mm_interconnect_0_sdram_s1_readdatavalid),                  //                                       .readdatavalid
		.sdram_s1_waitrequest                         (mm_interconnect_0_sdram_s1_waitrequest),                    //                                       .waitrequest
		.sdram_s1_chipselect                          (mm_interconnect_0_sdram_s1_chipselect),                     //                                       .chipselect
		.spi_ADC_spi_control_port_address             (mm_interconnect_0_spi_adc_spi_control_port_address),        //               spi_ADC_spi_control_port.address
		.spi_ADC_spi_control_port_write               (mm_interconnect_0_spi_adc_spi_control_port_write),          //                                       .write
		.spi_ADC_spi_control_port_read                (mm_interconnect_0_spi_adc_spi_control_port_read),           //                                       .read
		.spi_ADC_spi_control_port_readdata            (mm_interconnect_0_spi_adc_spi_control_port_readdata),       //                                       .readdata
		.spi_ADC_spi_control_port_writedata           (mm_interconnect_0_spi_adc_spi_control_port_writedata),      //                                       .writedata
		.spi_ADC_spi_control_port_chipselect          (mm_interconnect_0_spi_adc_spi_control_port_chipselect),     //                                       .chipselect
		.spi_DAC_spi_control_port_address             (mm_interconnect_0_spi_dac_spi_control_port_address),        //               spi_DAC_spi_control_port.address
		.spi_DAC_spi_control_port_write               (mm_interconnect_0_spi_dac_spi_control_port_write),          //                                       .write
		.spi_DAC_spi_control_port_read                (mm_interconnect_0_spi_dac_spi_control_port_read),           //                                       .read
		.spi_DAC_spi_control_port_readdata            (mm_interconnect_0_spi_dac_spi_control_port_readdata),       //                                       .readdata
		.spi_DAC_spi_control_port_writedata           (mm_interconnect_0_spi_dac_spi_control_port_writedata),      //                                       .writedata
		.spi_DAC_spi_control_port_chipselect          (mm_interconnect_0_spi_dac_spi_control_port_chipselect),     //                                       .chipselect
		.sync_in_s1_address                           (mm_interconnect_0_sync_in_s1_address),                      //                             sync_in_s1.address
		.sync_in_s1_write                             (mm_interconnect_0_sync_in_s1_write),                        //                                       .write
		.sync_in_s1_readdata                          (mm_interconnect_0_sync_in_s1_readdata),                     //                                       .readdata
		.sync_in_s1_writedata                         (mm_interconnect_0_sync_in_s1_writedata),                    //                                       .writedata
		.sync_in_s1_chipselect                        (mm_interconnect_0_sync_in_s1_chipselect),                   //                                       .chipselect
		.sysid_control_slave_address                  (mm_interconnect_0_sysid_control_slave_address),             //                    sysid_control_slave.address
		.sysid_control_slave_readdata                 (mm_interconnect_0_sysid_control_slave_readdata),            //                                       .readdata
		.uart_s1_address                              (mm_interconnect_0_uart_s1_address),                         //                                uart_s1.address
		.uart_s1_write                                (mm_interconnect_0_uart_s1_write),                           //                                       .write
		.uart_s1_read                                 (mm_interconnect_0_uart_s1_read),                            //                                       .read
		.uart_s1_readdata                             (mm_interconnect_0_uart_s1_readdata),                        //                                       .readdata
		.uart_s1_writedata                            (mm_interconnect_0_uart_s1_writedata),                       //                                       .writedata
		.uart_s1_begintransfer                        (mm_interconnect_0_uart_s1_begintransfer),                   //                                       .begintransfer
		.uart_s1_chipselect                           (mm_interconnect_0_uart_s1_chipselect),                      //                                       .chipselect
		.uart_dbg_s1_address                          (mm_interconnect_0_uart_dbg_s1_address),                     //                            uart_dbg_s1.address
		.uart_dbg_s1_write                            (mm_interconnect_0_uart_dbg_s1_write),                       //                                       .write
		.uart_dbg_s1_read                             (mm_interconnect_0_uart_dbg_s1_read),                        //                                       .read
		.uart_dbg_s1_readdata                         (mm_interconnect_0_uart_dbg_s1_readdata),                    //                                       .readdata
		.uart_dbg_s1_writedata                        (mm_interconnect_0_uart_dbg_s1_writedata),                   //                                       .writedata
		.uart_dbg_s1_begintransfer                    (mm_interconnect_0_uart_dbg_s1_begintransfer),               //                                       .begintransfer
		.uart_dbg_s1_chipselect                       (mm_interconnect_0_uart_dbg_s1_chipselect),                  //                                       .chipselect
		.VarSet_1_avalon_slave_address                (mm_interconnect_0_varset_1_avalon_slave_address),           //                  VarSet_1_avalon_slave.address
		.VarSet_1_avalon_slave_write                  (mm_interconnect_0_varset_1_avalon_slave_write),             //                                       .write
		.VarSet_1_avalon_slave_readdata               (mm_interconnect_0_varset_1_avalon_slave_readdata),          //                                       .readdata
		.VarSet_1_avalon_slave_writedata              (mm_interconnect_0_varset_1_avalon_slave_writedata),         //                                       .writedata
		.VarSet_1_avalon_slave_chipselect             (mm_interconnect_0_varset_1_avalon_slave_chipselect)         //                                       .chipselect
	);

	CPU_irq_mapper irq_mapper (
		.clk           (clk_clk),                            //       clk.clk
		.reset         (rst_controller_001_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),           // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),           // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),           // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),           // receiver3.irq
		.receiver4_irq (irq_mapper_receiver4_irq),           // receiver4.irq
		.receiver5_irq (irq_mapper_receiver5_irq),           // receiver5.irq
		.receiver6_irq (irq_mapper_receiver6_irq),           // receiver6.irq
		.sender_irq    (nios2_irq_irq)                       //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.reset_in1      (nios2_debug_reset_request_reset),    // reset_in1.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.clk            (clk_clk),                                //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_001_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_in1      (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

endmodule
